module top (
    // input
        input logic [7:0] data_i [1:0] ,
        input logic       clk_i        ,
        input logic       EA_i         ,
        input logic       EB_i         ,

    // output
        output logic [15:0] P_o 
     
);
    ex3 ex03(
        .*
    );

endmodule : top
