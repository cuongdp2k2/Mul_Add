module top (
    // input
        input logic  [7:0]   A_i        ,
        input logic          clk_i      ,

    // output
        output logic         overflow_o ,
                             carry_o    ,
        output logic [7:0]   S_o    
     
);
    main ex1(
        .*
    );

endmodule : top
